
//-----------------------------------------------------------------------------------------------------
//                                        VLSI Design Laboratory
//                               Istituto Nazionale di Fisica Nucleare (INFN)
//                                   via Giuria 1 10125, Torino, Italy
//-----------------------------------------------------------------------------------------------------
// [Filename]	    JTAG_MACRO.sv [RTL]
// [Project]	    RD53A pixel ASIC demonstrator
// [Author]         Luca Pacher - pacher@to.infn.it
// [Language]	    SystemVerilog 2012 [IEEE Std. 1800-2012]
// [Created]	    Jul  4, 2016
// [Modified]	    Jul 12, 2017
// [Description]    Top-level structural/RTL wrapper for the JTAG macro
// [Notes]          -
// [Status]         devel
//-----------------------------------------------------------------------------------------------------


// Dependencies:
//
// $RTL_DIR/eoc/jtag/JTAG_INSTRUCTION_REGISTER_codes_pkg.sv"
// $RTL_DIR/eoc/jtag/JTAG_TAP_FSM_codes_pkg.sv"
// $RTL_DIR/eoc/jtag/JTAG_TAP_FSM.sv
// $RTL_DIR/eoc/jtag/JTAG_INSTRUCTION_REGISTER.sv
// $RTL_DIR/eoc/jtag/JTAG_INSTRUCTION_DECODER.sv
// $RTL_DIR/eoc/jtag/JTAG_BYPASS_REGISTER.sv
// $RTL_DIR/eoc/jtag/JTAG_RX_REGISTER.sv
// $RTL_DIR/eoc/jtag/JTAG_TX_REGISTER.sv
// $RTL_DIR/eoc/jtag/JTAG_COMMAND_PULSER.sv
// $RTL_DIR/eoc/jtag/JTAG_AZ_REGISTER.sv
// $RTL_DIR/eoc/jtag/JTAG_AZ_GENERATOR.sv


`ifndef JTAG_MACRO__SV
`define JTAG_MACRO__SV


`timescale 1ns / 1ps
//`include "timescale.v"


`include "eoc/jtag/JTAG_INSTRUCTION_REGISTER_codes_pkg.sv"
`include "eoc/jtag/JTAG_TAP_FSM_codes_pkg.sv"
`include "eoc/jtag/JTAG_TAP_FSM.sv"
`include "eoc/jtag/JTAG_INSTRUCTION_REGISTER.sv"
`include "eoc/jtag/JTAG_INSTRUCTION_DECODER.sv"
`include "eoc/jtag/JTAG_BYPASS_REGISTER.sv"
`include "eoc/jtag/JTAG_RX_REGISTER.sv"
`include "eoc/jtag/JTAG_TX_REGISTER.sv"
`include "eoc/jtag/JTAG_COMMAND_PULSER.sv"
`include "eoc/jtag/JTAG_AZ_REGISTER.sv"
`include "eoc/jtag/JTAG_AZ_GENERATOR.sv"


module JTAG_MACRO (

   // standard JTAG I/O interface
   input  wire  JtagTrstB,                             // Test Reset (asynchronous, active low)      - from input PAD
   input  wire  JtagTck,                               // Test Clock                                 - from input PAD
   input  wire  JtagTms,                               // Test Mode Select                           - from input PAD
   input  wire  JtagTdi,                               // Test Data Input, sampled at posedge TCK    - from input PAD
   output logic JtagTdo,                               // Test Data Output, sampled at negedge TCK   - to tri-state output PAD

   output wire  JtagTdoEnable,                         // control signal for TDO tri-state output PAD
   output wire  JtagTapResetB,                         // optionally, feed the reset generated by TAP controller to user logic (TBD)


   // SER and DAC boundary scan chains
   output wire  JtagBoundaryScanShiftEn,
   output wire  JtagShiftDR,
   output wire  JtagUpdateDR,

   output wire  JtagBoundaryScanSerSel,                // select SER Boundary Scan Register (BSR)
   output wire  JtagBoundaryScanSerMode,               // control signal for SER BSC output multiplexer
   input  wire  JtagBoundaryScanSerTdo,                // serial data from SER BSR

   output wire  JtagBoundaryScanDacSel,                // select DAC Boundary Scan Register (BSR)
   output wire  JtagBoundaryScanDacMode,               // control signal for DAC BSC output multiplexer
   input  wire  JtagBoundaryScanDacTdo,                // serial data from DAC BSR


   // output data from JTAG ADDRESS register to bypass command-decoder FSM outputs [3:0] ChipID and [8:0] RegAddr
   output wire [3:0] JtagChipID,
   output wire [8:0] JtagRegAddr,


   // output data from JTAG CONFIGURATION register to bypass command-decoder FSM outputs [15:0] RegData
   output wire [15:0] JtagRegData,


   // output data from JTAG CALIBRATION register to bypass command-decoder FSM outputs [2:0] EdgeDelay, [5:0] EdgeWidth, [4:0] AuxDly, EdgeMode and AuxMode 
   output wire [2:0] JtagEdgeDly, 
   output wire [5:0] JtagEdgeWidth,
   output wire [4:0] JtagAuxDly,
   output wire       JtagEdgeMode,
   output wire       JtagAuxMode,


   // configuration data from JTAG GLOBALPULSE register to bypass command-decoder FSM ouputs [3:0] GlobalPulseWidth
   output wire [3:0] JtagGlobalPulseWidth,


   // single-pulse command flags to bypass command-decoder FSM outputs ECR, BCR, WrReg, RdReg, GenGlobalPulse and GenCal
   output wire JtagECR,
   output wire JtagBCR,
   output wire JtagWrReg,
   output wire JtagRdReg,
   output wire JtagGenGlobalPulse,
   output wire JtagGenCal,


   // 12-bit monitoring data + valid bit from ADC
   input  wire [12:0] JtagAdcData,


   // 128-bit readback data for READBACK register
   input  wire [127:0] JtagReadbackData,


   // PWM signal for Torino-only autozeroing
   output wire JtagPhiAZ,


   // nominal 160 MHz system clock
   input  wire Clk160, 


   // internal scan-chain interface (accessible through INSCAN instruction)
   output wire JtagInternalScanTdi,                                          // scan-in
   output wire JtagInternalScanEn,                                           // scan-en
   output wire JtagInternalScanMode,                                         // scan-mode
   input  wire JtagInternalScanTdo                                           // scan-out

   ) ;


   `ifndef ABSTRACT


   // some internal wires for interconnections

   wire TRST, TCK, TMS, TDI ;
   logic TDO ;

   wire SHIFT_DR, UPDATE_DR, CAPTURE_DR, CLOCK_DR ;
   wire SHIFT_IR, UPDATE_IR, CAPTURE_IR ;
   wire SELECT, ENABLE, TAP_RESET ;

   assign TRST = JtagTrstB ;
   assign TCK  = JtagTck   ;
   assign TMS  = JtagTms   ;
   assign TDI  = JtagTdi   ;

   assign JtagTdo       = TDO       ;
   assign JtagTdoEnable = ENABLE    ;
   assign JtagTapResetB = TAP_RESET ;
   assign JtagShiftDR   = SHIFT_DR  ;
   assign JtagUpdateDR  = UPDATE_DR ;

   wire TDO_BOUNDARYSCAN_SER, TDO_BOUNDARYSCAN_DAC ;

   assign TDO_BOUNDARYSCAN_SER = JtagBoundaryScanSerTdo ;
   assign TDO_BOUNDARYSCAN_DAC = JtagBoundaryScanDacTdo ;

   assign JtagBoundaryScanShiftEn = CLOCK_DR ;

   //-----------------------------------   TEST ACCESS PORT (TAP) CONTROLLER  ----------------------------------//

   JTAG_TAP_FSM  TAP (

      .TRST        (       TRST ),
      .TCK         (        TCK ),
      .TMS         (        TMS ),

      .SELECT_DR   (            ),
      .SHIFT_DR    (   SHIFT_DR ),
      .UPDATE_DR   (  UPDATE_DR ),
      .CAPTURE_DR  ( CAPTURE_DR ),
      .CLOCK_DR    (   CLOCK_DR ),           // **NOTE: used to enable shifting in boundary-scan registers

      .SELECT_IR   (            ),
      .SHIFT_IR    (   SHIFT_IR ),
      .UPDATE_IR   (  UPDATE_IR ),
      .CAPTURE_IR  ( CAPTURE_IR ),

      .RESET       (  TAP_RESET ),
      .SELECT      (     SELECT ),
      .ENABLE      (     ENABLE )

      ) ;



   //-----------------------------------------   INSTRUCTION REGISTER  -----------------------------------------//
 
   wire [4:0] OPCODE ;       // 5-bit JTAG instruction
   wire  TDO_IR ;            // TDO serial output from Instruction Register
   
   JTAG_INSTRUCTION_REGISTER  #( .DATA_WIDTH(5) ) INSTRUCTION_REGISTER (

      .RESET       ( /* TRST & */ TAP_RESET ),
      .CLOCK_IR    (                    TCK ),
      .SHIFT_IR    (               SHIFT_IR ),
      .CAPTURE_IR  (             CAPTURE_IR ),
      .UPDATE_IR   (              UPDATE_IR ),
      .TDI         (                    TDI ),
      .TDO         (                 TDO_IR ),
      .OPCODE      (            OPCODE[4:0] )

      ) ;




   //----------------------------------------   INSTRUCTION DECODER  -------------------------------------------//

   // selection flags for JTAG registers
   wire        ADDRESS_sel ;
   wire  CONFIGURATION_sel ;
   wire    CALIBRATION_sel ;
   wire    GLOBALPULSE_sel ;
   wire         BYPASS_sel ;
   wire         INSCAN_sel ;
   wire    AUTOZEROING_sel ;
   wire        ADCDATA_sel ;
   wire       READBACK_sel ;


   // command flags
   wire           WRREG_cmd ;
   wire           RDREG_cmd ;
   wire             ECR_cmd ;
   wire             BCR_cmd ;
   wire  GENGLOBALPULSE_cmd ;
   wire          GENCAL_cmd ;
   wire         STARTAZ_cmd ;
   wire          STOPAZ_cmd ;      


   JTAG_INSTRUCTION_DECODER  INSTRUCTION_DECODER (

      .OPCODE                (           OPCODE[4:0] ),
      .TCK                   (                   TCK ),
      .ADDRESS_sel           (           ADDRESS_sel ),
      .CONFIGURATION_sel     (     CONFIGURATION_sel ),
      .CALIBRATION_sel       (       CALIBRATION_sel ),
      .GLOBALPULSE_sel       (       GLOBALPULSE_sel ),
      .READBACK_sel          (          READBACK_sel ),
      .ADCDATA_sel           (           ADCDATA_sel ),
      .BYPASS_sel            (            BYPASS_sel ),
      .BOUNDARYSCAN_SER_sel  (  BOUNDARYSCAN_SER_sel ),
      .BOUNDARYSCAN_SER_mode ( BOUNDARYSCAN_SER_mode ),
      .BOUNDARYSCAN_DAC_sel  (  BOUNDARYSCAN_DAC_sel ),
      .BOUNDARYSCAN_DAC_mode ( BOUNDARYSCAN_DAC_mode ),
      .INSCAN_sel            (            INSCAN_sel ),
      .WRREG_cmd             (             WRREG_cmd ),
      .RDREG_cmd             (             RDREG_cmd ),
      .ECR_cmd               (               ECR_cmd ),
      .BCR_cmd               (               BCR_cmd ),
      .GENGLOBALPULSE_cmd    (    GENGLOBALPULSE_cmd ),
      .GENCAL_cmd            (            GENCAL_cmd ),
      .AUTOZEROING_sel       (       AUTOZEROING_sel ),
      .STARTAZ_cmd           (           STARTAZ_cmd ),
      .STOPAZ_cmd            (            STOPAZ_cmd )

      ) ;


   assign JtagBoundaryScanSerSel  = BOUNDARYSCAN_SER_sel ;
   assign JtagBoundaryScanSerMode = BOUNDARYSCAN_SER_mode ;

   assign JtagBoundaryScanDacSel  = BOUNDARYSCAN_DAC_sel ;
   assign JtagBoundaryScanDacMode = BOUNDARYSCAN_DAC_mode ;



   //------------------------------------------   BYPASS REGISTER  ---------------------------------------------//

   wire TDO_BYPASS ;

   JTAG_BYPASS_REGISTER   BYPASS_REGISTER (

      .CLOCK_DR   (                     TCK ),
      .SHIFT_DR   (   SHIFT_DR & BYPASS_sel ),
      .CAPTURE_DR ( CAPTURE_DR & BYPASS_sel ),
      .TDI        (                     TDI ),
      .TDO        (              TDO_BYPASS )

      ) ;



   //----------------------------------------   USER DATA REGISTERS  -------------------------------------------//


   // 14-bit ADDRESS register, bypass [8:0] RegAddr and [3:0] ChipID outputs from command-decoder FSM and set the normal/autoincrement mode

   wire TDO_ADDRESS ;
   wire [13:0] ADDRESS_reg ;
 
   JTAG_RX_REGISTER   #( .DATA_WIDTH(14) ) ADDRESS_REGISTER (

      .RESET      (  /* TRST & */ TAP_RESET ),
      .CLOCK_DR   (                     TCK ),
      .SHIFT_DR   (  SHIFT_DR & ADDRESS_sel ),
      .UPDATE_DR  ( UPDATE_DR & ADDRESS_sel ),
      .TDI        (                     TDI ),
      .TDO        (             TDO_ADDRESS ),
      .SHADOW     (       ADDRESS_reg[13:0] )

      ) ;

   assign JtagChipID   = ADDRESS_reg [ 3:0] ;
   assign JtagRegAddr  = ADDRESS_reg [12:4] ;

   wire   normal0_auto1 ;
   assign normal0_auto1 = ADDRESS_reg [13] ;


   // 16-bit CONFIGURATION register, bypass [15:0] RegData outputs from command-decoder FSM

   wire TDO_CONFIGURATION ;
   wire [15:0] CONFIGURATION_reg ;

   JTAG_RX_REGISTER   #( .DATA_WIDTH(16) ) CONFIGURATION_REGISTER (

      .RESET      (        /* TRST & */ TAP_RESET ),
      .CLOCK_DR   (                           TCK ),
      .SHIFT_DR   (  SHIFT_DR & CONFIGURATION_sel ),
      .UPDATE_DR  ( UPDATE_DR & CONFIGURATION_sel ),
      .TDI        (                           TDI ),
      .TDO        (             TDO_CONFIGURATION ),
      .SHADOW     (       CONFIGURATION_reg[15:0] )

      ) ;

   assign JtagRegData = CONFIGURATION_reg ;



   // 16-bit CALIBRATION register, bypass [2:0] EdgeDly, [5:0] EdgeWidth, [4:0] AuxDly, EdgeMode and AuxMode outputs from command-decoder FSM

   wire TDO_CALIBRATION ;
   wire [15:0] CALIBRATION_reg ;

   JTAG_RX_REGISTER   #( .DATA_WIDTH(16) ) CALIBRATION_REGISTER (

      .RESET      (      /* TRST */ & TAP_RESET ),
      .CLOCK_DR   (                         TCK ),
      .SHIFT_DR   (  SHIFT_DR & CALIBRATION_sel ),
      .UPDATE_DR  ( UPDATE_DR & CALIBRATION_sel ),
      .TDI        (                         TDI ),
      .TDO        (             TDO_CALIBRATION ),
      .SHADOW     (       CALIBRATION_reg[15:0] )

      ) ;

   assign JtagEdgeDly   = CALIBRATION_reg [ 2:0] ;
   assign JtagEdgeWidth = CALIBRATION_reg [ 8:3] ;
   assign JtagAuxDly    = CALIBRATION_reg [13:9] ;
   assign JtagEdgeMode  = CALIBRATION_reg [14  ] ;
   assign JtagAuxMode   = CALIBRATION_reg [15  ] ;



   // 4-bit GLOBALPULSE register, bypass [3:0] GlobalPulseWidth outputs from command-decoder FSM

   wire TDO_GLOBALPULSE ;
   wire [3:0] GLOBALPULSE_reg ;

   JTAG_RX_REGISTER   #( .DATA_WIDTH(4) ) GLOBALPULSE_REGISTER (

      .RESET      (      /* TRST & */ TAP_RESET ),
      .CLOCK_DR   (                         TCK ),
      .SHIFT_DR   (  SHIFT_DR & GLOBALPULSE_sel ),
      .UPDATE_DR  ( UPDATE_DR & GLOBALPULSE_sel ),
      .TDI        (                         TDI ),
      .TDO        (             TDO_GLOBALPULSE ),
      .SHADOW     (        GLOBALPULSE_reg[3:0] )

      ) ;

   assign JtagGlobalPulseWidth = GLOBALPULSE_reg ;




   // 13-bit readout register for monitoring data from ADC

   wire TDO_ADCDATA ;

   JTAG_TX_REGISTER   #( .DATA_WIDTH(13) ) ADC_REGISTER (

      .RESET      (   /* TRST & */ TAP_RESET ),
      .CLOCK_DR   (                      TCK ),
      .CAPTURE_DR ( CAPTURE_DR & ADCDATA_sel ),
      .SHIFT_DR   (   SHIFT_DR & ADCDATA_sel ),
      .PDATA      (        JtagAdcData[12:0] ),
      .TDI        (                      TDI ),
      .TDO        (              TDO_ADCDATA )

      ) ;



   // 128-bit readout register for readback data from DCB

   wire TDO_READBACK ;

   JTAG_TX_REGISTER   #( .DATA_WIDTH(128) ) READBACK_REGISTER (

      .RESET      (    /* TRST & */ TAP_RESET ),
      .CLOCK_DR   (                       TCK ),
      .CAPTURE_DR ( CAPTURE_DR & READBACK_sel ),
      .SHIFT_DR   (   SHIFT_DR & READBACK_sel ),
      .PDATA      (   JtagReadbackData[127:0] ),
      .TDI        (                       TDI ),
      .TDO        (              TDO_READBACK )

      ) ;



   // 27-bit Torino-only AUTOZEROING register

   wire TDO_AUTOZEROING ;
   wire [26:0] AUTOZEROING_reg ;

   JTAG_AZ_REGISTER  AUTOZEROING_REGISTER ( 

      .RESET      (        /* TRST &*/ TAP_RESET ),
      .CLOCK_DR   (                          TCK ),
      .CAPTURE_DR ( CAPTURE_DR & AUTOZEROING_sel ),
      .SHIFT_DR   (   SHIFT_DR & AUTOZEROING_sel ),
      .UPDATE_DR  (  UPDATE_DR & AUTOZEROING_sel ),
      .TDI        (                          TDI ),
      .TDO        (              TDO_AUTOZEROING ),
      .SHADOW     (        AUTOZEROING_reg[26:0] )

      ) ;



   //-----------------------------------   INTERNAL SCAN-CHAIN INTERFACE  --------------------------------------//

   
   assign JtagInternalScanMode = INSCAN_sel ;
   assign JtagInternalScanEn   = INSCAN_sel & SHIFT_DR ;

   wire   TDO_INSCAN ;
   assign TDO_INSCAN = JtagInternalScanTdo ;

   assign JtagInternalScanTdi = TDI & INSCAN_sel ;



   //-------------------------------------   TDO OUTPUT DECODING LOGIC  ----------------------------------------//


   // Data Registers (DR) multiplexing logic depending on Instruction Decoder outputs

   logic TDO_DR ;

   always_comb begin

      // TDO_DR = 1'b0 ;
      TDO_DR = TDO_BYPASS ;

      if( BYPASS_sel == 1'b1 )
         TDO_DR = TDO_BYPASS ;

      else if( BOUNDARYSCAN_SER_sel == 1'b1 )
         TDO_DR = TDO_BOUNDARYSCAN_SER ;

      else if( BOUNDARYSCAN_DAC_sel == 1'b1 )
         TDO_DR = TDO_BOUNDARYSCAN_DAC ;

      else if( INSCAN_sel == 1'b1 )
         TDO_DR = TDO_INSCAN ;

      else if( ADDRESS_sel == 1'b1 )
         TDO_DR = TDO_ADDRESS ;

      else if( CONFIGURATION_sel == 1'b1 )
         TDO_DR = TDO_CONFIGURATION ;

      else if( CALIBRATION_sel == 1'b1 )
         TDO_DR = TDO_CALIBRATION ;

      else if( GLOBALPULSE_sel == 1'b1 )
         TDO_DR = TDO_GLOBALPULSE ;

      else if( ADCDATA_sel == 1'b1 )
         TDO_DR = TDO_ADCDATA ;

      else if( READBACK_sel == 1'b1 )
         TDO_DR = TDO_READBACK ;

      else if( AUTOZEROING_sel == 1'b1 )
         TDO_DR = TDO_AUTOZEROING ;

      else 
         TDO_DR = TDO_BYPASS ;

   end  // always_comb




   // Data Registers/Instruction Register TDO multiplexer
   wire   TDO_mux ;
   assign TDO_mux = ( SELECT == 1'b1 ) ? TDO_IR : TDO_DR ;


   // output DFF
   always_ff @(negedge TCK) begin     // **NOTE: according to IEEE Std. 1149.1-2001, TDO must change at NEGATIVE edge of TCK (no reset is foreseen for this output DFF)
      TDO <= TDO_mux ;
   end



   //------------------------------------------   COMMAND PULSER  ----------------------------------------------//

   // automatically generate a WrReg flag from UPDATE_DR when in auto-increment mode

   logic WRREG_auto ;

   always_ff @(posedge TCK)
      WRREG_auto <= UPDATE_DR & CONFIGURATION_sel & normal0_auto1 ;


   JTAG_COMMAND_PULSER COMMAND_PULSER (

      .Clk160              (                 Clk160 ),
      .JtagTck             (                JtagTck ),
      .WRREG_cmd           ( WRREG_cmd | WRREG_auto ),
      .RDREG_cmd           (              RDREG_cmd ),
      .ECR_cmd             (                ECR_cmd ),
      .BCR_cmd             (                BCR_cmd ),
      .GENGLOBALPULSE_cmd  (     GENGLOBALPULSE_cmd ),
      .GENCAL_cmd          (             GENCAL_cmd ),
      .JtagWrReg           (              JtagWrReg ),
      .JtagRdReg           (              JtagRdReg ),
      .JtagECR             (                JtagECR ),
      .JtagBCR             (                JtagBCR ),
      .JtagGenGlobalPulse  (     JtagGenGlobalPulse ),
      .JtagGenCal          (             JtagGenCal )

      ) ;



   //------------------------------------   AUTOZEROING PWM GENERATOR  -----------------------------------------//


   wire [ 4:0] Ndelay ;
   wire [ 7:0] Nhigh ;
   wire [13:0] Nlow ;

   assign Ndelay = AUTOZEROING_reg[ 4: 0] ;
   assign Nhigh  = AUTOZEROING_reg[12: 5] ;
   assign Nlow   = AUTOZEROING_reg[26:13] ;


   JTAG_AZ_GENERATOR  AUTOZEROING_GENERATOR (

      .RESET       ( /*TRST & */ TAP_RESET ),
      .TCK         (                   TCK ),
      .STARTAZ     (           STARTAZ_cmd ),           
      .STOPAZ      (            STOPAZ_cmd ),
      .NDELAY      (           Ndelay[4:0] ), 
      .NHIGH       (            Nhigh[7:0] ),
      .NLOW        (            Nlow[13:0] ),
      .JTAG_PHI_AZ (             JtagPhiAZ )

      ) ;


   `endif   // ABSTRACT

endmodule : JTAG_MACRO

`endif   // JTAG_MACRO__SV


//-----------------------------------------------------------------------------------------------------
// [Filename]       Cmd.sv [RTL]
// [Project]        RD53A pixel ASIC demonstrator
// [Author]         Roberto Beccherle - Roberto.Beccherle@cern.ch
// [Language]       SystemVerilog 2012 [IEEE Std. 1800-2012]
// [Created]        Feb 03, 2017
// [Modified]       Feb 03, 2017
// [Description]    Command Decoder
// [Notes]          Reset is Synchronous and active low
//                  All signals generated by the Comand Decoder are active one clock cycle before the 40MHz clock is rising
//                  CalAux, CalEdge and GlobalPulse with delay = 0 start with the rising edge of the 40 MHz clock 
// [Version]        2.0
// [Status]         devel
//-----------------------------------------------------------------------------------------------------


// Dependencies:
//
// $RTL_DIR/eoc/cmd/Cmd_FSM.sv
// $RTL_DIR/eoc/cmd/GenCal.sv
// $RTL_DIR/eoc/cmd/GenGlobalPulse.sv
//-----------------------------------------------------------------------------------------------------


`ifndef CMD_SV 
`define CMD_SV

//#
//# Timescale directive
//`include "Timescale.v"
//# All definitions of signals relative to the Command Decoder
`include "eoc/cmd/Cmd_FSM.sv"
`include "eoc/cmd/GenCal.sv"
`include "eoc/cmd/GenGlobalPulse.sv"
// 
// Command Decoder FSM
// These are the commands supported and their format
// BCR:         {Bcr,Bcr} --> Generate BCR pulse
// ECR:         {Ecr,Ecr} --> Generate ECR pulse
// CAL:         {Cal,Cal}{ChipId[3:0],CalEdgeMode,CalEdgeDelay[2:0],CalEdgeWidth[5:4]}{CalEdgeWidth[3:0],CalAuxMode,CalAuxDly[4:0]}  [Cal +DD +DD] --> Genrate CalEdge, CalAux
//                                  0=step 1=pulse,1 to 8 @  40MHz , 0 to 63 @ 160MHz, 0 to 63 @ 160MHz ,  SetTo   ,1 to 32 @ 160MHz
// GlobalPulse: {GlobalPulse,GlobalPulse}{ChipId[3:0],0, GlobalPulseWidth[3:0],0} Generate GlobalPulse signal and GlobalPulseWidth bus. [widths are 1,2,4,8,16,32,64,128,256,512]
// WrReg: (0)   {WrReg,WrReg} {{ChipId[3:0],WrRegMode,Addr[8:4]} {Addr[3:0],Data[15:10]} {Data[9:0]} [WrReg +DD +DD +DD]
//  ...   (1)   {Data[15:6]} {Data[5:0],Data[15:12]} {Data[11:2]} {Data[1:0],Data[15:7]} {Data[6:0],Data[15:8]} {Data[7:0],Data[15:9]} {Data[8:0],Data[15:10]} {Data[9:0]} [+DD +DD +DD +DD +DD +DD +DD +DD]
// Rrdeg:       {RdReg,RdReg} {{ChipId[3:0],0,Addr[8:4]} {Addr[3:0],0_0000} {Data[9:0]} [RdReg +DD +DD]
// Null:        {Null, Null} No command, just ignore it
//-----------------------------------------------------------------------------------------------------
// In case of the chip goes out of sync (Sync = 1'b0) the command decoder will stop working, going back to SYNC state
//-----------------------------------------------------------------------------------------------------
// 
// 


module Cmd(
       //
       // Command Decoder 
       //
       // Outputs
       output logic        Trigger,        // Trigger signal
       output logic  [4:0] TriggerTag,     // The correct 7 bit tag
       output logic        ECR,            // Event Counter Reset
       output logic        CalEdge,        // Only if ChipId matches
       output logic        CalAux,         // Only if ChipId matches
       output logic        RdReg,          // Only if ChipId matches
       output logic        WrReg,          // Only if ChipId matches
       output logic        GlobalPulse,    // Only if ChipId matches
       output logic  [8:0] RegAddr,        // Address of the register
       output logic [15:0] RegData,        // Data to be written in the addressed register
       output wire  [15:0] BCIDCnt,        // BCID counter value
       output logic [15:0] TrigCnt,        // Trigger counter value
       output logic [15:0] ErrCnt,         // Error counter value
       output logic        CmdErr,         // There is an Error
       output logic [15:0] BitFlipWngCnt,  // BitFlip Warning  counter value
       output logic        BitFlipWng,     // There is a BitFlip warning
       output logic [15:0] BitFlipErrCnt,  // BitFlip Error counter value
       output logic        BitFlipErr,     // There is a BitFlip error
       // External Trigger signal coming from a Pad
       input  wire         ExtTrigger, // Is a pull down
       // Input signals coming from JTAG block, to be muxed inside the Command Decoder
       input  wire         BypassCmd,
       input  wire         JtagTck,
       input  wire [ 3:0]  JtagChipID,
       input  wire [ 8:0]  JtagRegAddr,
       input  wire [15:0]  JtagRegData,
       input  wire [ 2:0]  JtagEdgeDly,
       input  wire [ 5:0]  JtagEdgeWidth,
       input  wire [ 4:0]  JtagAuxDly,
       input  wire         JtagEdgeMode,
       input  wire         JtagAuxMode,
       input  wire [ 3:0]  JtagGlobalPulseWidth,
       input  wire         JtagWrReg,
       input  wire         JtagRdReg,
       input  wire         JtagECR,
       input  wire         JtagBCR,
       input  wire         JtagGenGlobalPulse,
       input  wire         JtagGenCal,
       // Inputs
       input  wire        clk, 
       input  wire        Reset_b,     // Synchronous active low
       input  wire         WrBCIDCnt,   // Resets the BCID Counter
       input  wire         WrTrigCnt,   // Resets the Trigger Counter
       input  wire   WrBitFlipWngCnt,   // Resets the Bit Flip Warning Counter
       input  wire   WrBitFlipErrCnt,   // Resets the Bit Flip Error Counter
       input  wire          WrErrCnt,   // Resets the Error Counter

       input  wire [15:0] Input,   // Input data (stable for 16 clk cycles)
       input  wire  [2:0] ChipId,  // ChipId coming from wire bnd pads
       input  wire        Locked,  // Input is locked, we expect data
       input  wire        Load     // Active when data is stable (1 clk cycle every 16)
       );


//
// Local signal definition
//
logic [15:0] TimCnt, CmdRegData, RegData_mux, InputFSM;
logic  [8:0] CmdRegAddr, RegAddr_mux;
logic  [5:0] EdgeWidth_mux, CmdEdgeWidth;
logic  [2:0] EdgeDly_mux, CmdEdgeDly;
logic  [4:0] AuxDly_mux, CmdAuxDly;
logic        EdgeMode_mux, CmdEdgeMode;
logic        AuxMode_mux, CmdAuxMode;
logic  [3:0] GlobalPulseWidth_mux, CmdGlobalPulseWidth;
logic  [3:0] ChipId_mux, CmdChipId;
logic  [4:0] TrgTagFsm;
logic        Trigger1, Trigger2, Trigger3, Trigger4, Trigger_comb, Trigger_mux,
             TrgFsm1, TrgFsm2, TrgFsm3, TrgFsm4,
             BCR_mux, CmdBCR, ECR_mux, CmdECR, 
             BitFlipWarning, BitFlipWarningFsm, BitFlipWarning_comb,
             Error, ErrorFsm, Error_comb,
             BitFlipError, BitFlipErrorFsm, BitFlipError_comb, 
             FSM_Reset_b,                           // Cmd_FSM reaset signal
             ChipIdOK,
             GenCal_mux, CmdGenCal, 
             GenGlobalPulse_mux, CmdGenGlobalPulse,
             GPDelay1, GPDelay2,                    // Used to align GlobalPulse signal
             RdReg_mux, CmdRdReg,  
             WrReg_mux, CmdWrReg, 
             CmdIncrBCID, 
             CmdBCIDCntRst,      // Reset the BCID counter
             TrigCntRst,         // Reset the Trigger counter
             ErrCntRst,          // Reset the Error counter
             BitFlipWngCntRst,   // Reset the Bit Flip Warning counter
             BitFlipErrCntRst;   // Reset the Bit Flip Error counter

// synopsys sync_set_reset "Reset_b"
             
//
//                    ###       ##       ##               ###
// ##   ##             ##       ##       ##                ##
// ##   ##             ##       ##                         ##
// ### ###  ##   ##    ##     ######   ####     ######     ##      #####   ##  ##    #####   ## ###    #####
// ## # ##  ##   ##    ##       ##       ##     ##   ##    ##     ##   ##   ####    ##   ##  ###      ##
// ## # ##  ##   ##    ##       ##       ##     ##   ##    ##     #######    ##     #######  ##        ####
// ##   ##  ##  ###    ##       ##       ##     ##   ##    ##     ##        ####    ##       ##           ##
// ##   ##   ### ##   ####       ###   ######   ######    ####     #####   ##  ##    #####   ##       #####
//                                              ##
//                                              ##
//
//
// Multiplexers between JTAG and Command Decoder FSM signals
//
assign ChipId_mux[3:0]            =  ( BypassCmd == 1'b1 )  ?  JtagChipID[3:0]           :  CmdChipId[3:0] ;
assign RegAddr_mux[8:0]           =  ( BypassCmd == 1'b1 )  ?  JtagRegAddr[8:0]          :  CmdRegAddr[8:0] ;
assign RegData_mux[15:0]          =  ( BypassCmd == 1'b1 )  ?  JtagRegData[15:0]         :  CmdRegData[15:0] ;
assign EdgeWidth_mux[5:0]         =  ( BypassCmd == 1'b1 )  ?  JtagEdgeWidth[5:0]        :  CmdEdgeWidth[5:0] ;
assign EdgeDly_mux[2:0]           =  ( BypassCmd == 1'b1 )  ?  JtagEdgeDly[2:0]          :  CmdEdgeDly[2:0] ;
assign AuxDly_mux[4:0]            =  ( BypassCmd == 1'b1 )  ?  JtagAuxDly[4:0]           :  CmdAuxDly[4:0] ;
assign EdgeMode_mux               =  ( BypassCmd == 1'b1 )  ?  JtagEdgeMode              :  CmdEdgeMode ;
assign AuxMode_mux                =  ( BypassCmd == 1'b1 )  ?  JtagAuxMode               :  CmdAuxMode ;
assign GenCal_mux                 =  ( BypassCmd == 1'b1 )  ?  JtagGenCal                :  CmdGenCal ;
assign GlobalPulseWidth_mux[3:0]  =  ( BypassCmd == 1'b1 )  ?  JtagGlobalPulseWidth[3:0] :  CmdGlobalPulseWidth[3:0] ;
assign GenGlobalPulse_mux         =  ( BypassCmd == 1'b1 )  ?  JtagGenGlobalPulse        :  CmdGenGlobalPulse ;


//
// BCR command
assign BCR_mux   =  ( BypassCmd == 1'b1 ) ? JtagBCR   : TimCnt[1] & CmdBCR;
//
// ECR command
assign ECR_mux   =  ( BypassCmd == 1'b1 ) ? JtagECR   : TimCnt[1] & CmdECR;
//
// RdReg command
assign RdReg_mux =  ( BypassCmd == 1'b1 ) ? JtagRdReg : TimCnt[1] & CmdRdReg & ChipIdOK;
//
// WrReg command
assign WrReg_mux =  ( BypassCmd == 1'b1 ) ? JtagWrReg : TimCnt[1] & CmdWrReg & ChipIdOK;

//
// Multiplexer for Trigger
assign Trigger_mux         = ( BypassCmd == 1'b1 ) ? ExtTrigger :  Trigger_comb  ; 

//
// Cmd_FSM reset signal: it is also reset when Locked is low (no lock on channel)
assign FSM_Reset_b = Reset_b & Locked; 

//
// Delayed GlobalPulse
assign GlobalPulse = GPDelay2;

//
// ChipIdOK is set when ChipIdFsm matches ChipId, or we are in broadcast
assign ChipIdOK     = ChipId_mux[3] | (ChipId_mux[2:0] == ChipId[2:0]);
//
// Trigger 
assign        Trigger1 = TimCnt[1]  & TrgFsm1;
assign        Trigger2 = TimCnt[5]  & TrgFsm2;
assign        Trigger3 = TimCnt[9]  & TrgFsm3;
assign        Trigger4 = TimCnt[13] & TrgFsm4;
assign    Trigger_comb = Trigger1 | Trigger2 | Trigger3 | Trigger4;
//
// Trigger Tag
assign TriggerTag = TrgTagFsm;
//
// Increment the BCID counter each time there is a 40 MHz clock
assign CmdIncrBCID = TimCnt[2] | TimCnt[6] | TimCnt[10] | TimCnt[14] ;
//
// Trigger counter is incremented each time there is a Trigger
// and cleared by a reset, an ECR or a WrTrigCnt
assign TrigCntRst = (Reset_b == 1'b0) | ECR | WrTrigCnt;
//
// BitFlip Warning signal
assign BitFlipWarning_comb = TimCnt[0] & BitFlipWarningFsm;
//
// BitFlip Error signal
assign BitFlipError_comb   = TimCnt[0] & BitFlipErrorFsm;
//
// Error signal
assign Error_comb   = TimCnt[0] & ErrorFsm;
//
// Signal to sample next_state transition (has to be one clk cycle after Load)
logic  Sample;
assign Sample = TimCnt[0];
//
// Counter Reset signals
//
assign    CmdBCIDCntRst = (Reset_b == 1'b0) | BCR_mux | WrBCIDCnt;  // Cleared by a reset, a BCR or a WrReg command
assign BitFlipWngCntRst = (Reset_b == 1'b0) | WrBitFlipWngCnt;      // Cleared by a reset or a WrReg command
assign BitFlipErrCntRst = (Reset_b == 1'b0) | WrBitFlipErrCnt;      // Cleared by a reset or a WrReg command
assign        ErrCntRst = (Reset_b == 1'b0) | WrErrCnt;             // Cleared by a reset or a WrReg command



//
//                        ##            ###
// ##   ##                ##             ##
// ##   ##                ##             ##
// ### ###   #####    ######  ##   ##    ##      #####    #####
// ## # ##  ##   ##  ##   ##  ##   ##    ##     ##   ##  ##
// ## # ##  ##   ##  ##   ##  ##   ##    ##     #######   ####
// ##   ##  ##   ##  ##   ##  ##  ###    ##     ##           ##
// ##   ##   #####    ######   ### ##   ####     #####   #####
//
//
//
//
// Instantiate the Command Decoder FSM
Cmd_FSM  Cmd_FSM_i (

   // Inputs
   .clk              (                      clk ),
   .Reset_b          (              FSM_Reset_b ),
   .Input            (           InputFSM[15:0] ),
   .Enable           (                     Load ),
   .Sample           (                   Sample ),

   // Outputs are all registered
   .Trigger1         (                  TrgFsm1 ),
   .Trigger2         (                  TrgFsm2 ),
   .Trigger3         (                  TrgFsm3 ),
   .Trigger4         (                  TrgFsm4 ),
   .TriggerTag       (                TrgTagFsm ),
   .ECR              (                   CmdECR ),
   .BCR              (                   CmdBCR ),
   .RdReg            (                 CmdRdReg ),
   .WrReg            (                 CmdWrReg ), 
   .RegData          (         CmdRegData[15:0] ),
   .RegAddr          (          CmdRegAddr[8:0] ),
   .ChipId           (           CmdChipId[3:0] ),
   .GlobalPulseWidth ( CmdGlobalPulseWidth[3:0] ),
   .GenGlobalPulse   (        CmdGenGlobalPulse ),
   .EdgeWidth        (        CmdEdgeWidth[5:0] ),
   .EdgeDly          (          CmdEdgeDly[2:0] ),
   .AuxDly           (           CmdAuxDly[4:0] ),
   .EdgeMode         (              CmdEdgeMode ),
   .AuxMode          (               CmdAuxMode ),
   .GenCal           (                CmdGenCal ),
   .BitFlipWarning   (        BitFlipWarningFsm ),     // True if there has been a BitFlip and it has been corrected
   .BitFlipError     (          BitFlipErrorFsm ),     // True if there has been a Bit Flip in any Symbol (and it has not been corrected)
   .Error            (                 ErrorFsm )      // True if nothing matched in SYNC or DATA states or if a Command Counter has a wrong vaulue

   ) ;

// 
// Instantiate the Calibration pulse generator 

GenCal  GenCal_i (

   // Inputs
   .clk       (                   clk ), 
   .Reset_b   (               Reset_b ),      // Syncronous reset active low
   .EdgeWidth (    EdgeWidth_mux[5:0] ),      // from 0 to 63
   .EdgeDly   (      EdgeDly_mux[2:0] ),      // from 1 to 8
   .AuxDly    (       AuxDly_mux[4:0] ),      // from 1 to 32
   .GenCal    ( GenCal_mux & ChipIdOK ),      // Generate Cal pulses only if ChipId matches
   .EdgeMode  (          EdgeMode_mux ),      // Step (EdgeMode = 0) or Pulse (EdgeMode = 1)
   .AuxMode   (           AuxMode_mux ),      // Determines the value of the aux signal

    // Outputs [Are all registered]
    .CalEdge  (               CalEdge ), 
    .CalAux   (                CalAux )

   ) ;

// 
// Instantiate the Calibration pulse generator

wire GlobalPulse_int ;
 
GenGlobalPulse  GenGlobalPulse_i (

   // Inputs
  .clk              (                           clk ),
  .Reset_b          (                       Reset_b ), // Syncronous reset active low
  .GlobalPulseWidth (     GlobalPulseWidth_mux[3:0] ),
  .GenGlobalPulse   ( GenGlobalPulse_mux & ChipIdOK ), // Generate GlobalPulse only if ChipId matches

   // Outputs
   .GlobalPulse     (               GlobalPulse_int )

   ) ;

// 
// Shift Register to generate timing of signals
// Each time there is a Load we write 16'b1 to the SR
always_ff @(posedge clk) begin: TimingCounter
    if (Reset_b == 1'b0) TimCnt <=   'b0;
    else if (Load)       TimCnt <= 16'b1;
    else                 TimCnt <= {TimCnt[14:0],1'b0};
end: TimingCounter

// //
// // Set Trigger specific Tags
// always_ff @(posedge clk) begin : proc_TrgTag
//     if (Load == 1'b1) begin 
//         TriggerTag[6:5] <= 'b0;
//     end else begin
//         if(Trigger1) TriggerTag[6:5] <= 2'b00;
//         if(Trigger2) TriggerTag[6:5] <= 2'b01;
//         if(Trigger3) TriggerTag[6:5] <= 2'b10;
//         if(Trigger4) TriggerTag[6:5] <= 2'b11;
//     end // end else
// end // proc_TrgTag

// 
// Register all Outputs
always_ff @(posedge clk) begin: RegOutputs_AFF
    if (Reset_b == 1'b0) begin
        BitFlipWarning <= 'b0;
        BitFlipError   <= 'b0;
        Error          <= 'b0;
        Trigger        <= 'b0;
        ECR            <= 'b0;
        RdReg          <= 'b0;
        WrReg          <= 'b0;
        RegAddr        <= 'b0;
        RegData        <= 'b0;
        GPDelay1       <= 'b0;
        GPDelay2       <= 'b0;
    end else begin
        BitFlipWarning <= BitFlipWarning_comb;
        BitFlipError   <= BitFlipError_comb;
        Error          <= Error_comb;
        Trigger        <= Trigger_mux;
        ECR            <= ECR_mux;
        RdReg          <= RdReg_mux;
        WrReg          <= WrReg_mux;
        RegAddr        <= RegAddr_mux;
        RegData        <= RegData_mux;
        GPDelay1       <= GlobalPulse_int;
        GPDelay2       <= GPDelay1;
    end
end: RegOutputs_AFF

always_ff @(posedge clk) begin : proc_dlyinput
    InputFSM     <= Input;
end // proc_dlyinput

// 
// Counter to keep track of the Bunch Crossing

logic [15:0] CmdBCIDCnt ; 

always_ff @(posedge clk) begin: CmdBCIDCounter
    if (CmdBCIDCntRst == 1'b1)
       CmdBCIDCnt <= 'b0;
    else if (CmdIncrBCID)
       CmdBCIDCnt <= CmdBCIDCnt + 1;
    else
       CmdBCIDCnt <= CmdBCIDCnt;
end: CmdBCIDCounter


//////////////////////////////////////////////
//   **BACKUP: BCID counter from JTAG       //
//////////////////////////////////////////////

// clock gating
logic BypassCmd_latch ;

always_latch begin
   if( JtagTck == 1'b0 )
      BypassCmd_latch <= BypassCmd ;
end 


wire JtagTck_gated ;
assign JtagTck_gated = JtagTck & BypassCmd_latch ;

// BCID counter using JTAG TCK

wire JtagBCIDCntRst = (Reset_b == 1'b0) | JtagBCR ;

logic [15:0] JtagBCIDCnt ;

always_ff @(posedge JtagTck_gated ) begin : JtagBCIDCounter

   if( JtagBCIDCntRst == 1'b1 )
      JtagBCIDCnt <= 'b0 ;

   else
      JtagBCIDCnt <= JtagBCIDCnt + 1 ;

end : JtagBCIDCounter


assign BCIDCnt = ( BypassCmd == 1'b1 ) ? JtagBCIDCnt : CmdBCIDCnt ; 


// 
// Counter to keep track of Triggers
always_ff @(posedge clk) begin: TrigCounter
    if (TrigCntRst == 1'b1) TrigCnt <= 'b0;
    else if (Trigger)       TrigCnt <= TrigCnt + 1;
    else                    TrigCnt <= TrigCnt;
end: TrigCounter

// 
// Counter to keep track of Errors
always_ff @(posedge clk) begin: ErrorCounter
    if (ErrCntRst == 1'b1) ErrCnt <= 'b0;
    else if (Error)        ErrCnt <= ErrCnt + 1;
    else                   ErrCnt <= ErrCnt;
end: ErrorCounter 

//
// CmdErr generator
always_ff @(posedge clk) begin: CmdErrGenerator
    if (ErrCnt == 16'b0) CmdErr <= 1'b0;
    else                 CmdErr <= 1'b1;
end: CmdErrGenerator

// 
// Counter to keep track of BitFlip warnings
always_ff @(posedge clk) begin: BitFlipWngCounter
    if (BitFlipWngCntRst == 1'b1) BitFlipWngCnt <= 'b0;
    else if (BitFlipWarning)      BitFlipWngCnt <= BitFlipWngCnt + 1;
    else                          BitFlipWngCnt <= BitFlipWngCnt;
end: BitFlipWngCounter

//
// BitFlipWng generator
always_ff @(posedge clk) begin: BitFlipWngGenerator
    if (BitFlipWngCnt == 16'b0) BitFlipWng <= 1'b0;
    else                        BitFlipWng <= 1'b1;
end: BitFlipWngGenerator

// 
// Counter to keep track of BitFlip errors
always_ff @(posedge clk) begin: BitFlipErrCounter
    if (BitFlipErrCntRst == 1'b1) BitFlipErrCnt <= 'b0;
    else if (BitFlipError)        BitFlipErrCnt <= BitFlipErrCnt + 1;
    else                          BitFlipErrCnt <= BitFlipErrCnt;
end: BitFlipErrCounter

//
// BitFlipErr generator
always_ff @(posedge clk) begin: BitFlipErrGenerator
    if (BitFlipErrCnt == 16'b0) BitFlipErr <= 1'b0;
    else                        BitFlipErr <= 1'b1;
end: BitFlipErrGenerator

endmodule : Cmd

`endif // CMD_SV

// Library - RD53_IO, Cell - RD53_TOP_BLOCKS, View - schematic
// LAST TIME SAVED: Jun 28 15:51:55 2017
// NETLIST TIME: Jun 29 14:52:06 2017

module RD53_TOP_BLOCKS ( BGPV_OE12, BGPV_OE34, BGPV_OE56, BGPV_PA1,
     BGPV_PA2, BGPV_PA3, BGPV_PA4, BGPV_PA5, BGPV_PA6, BGPV_SF_IN,
     BGPV_SF_OUT, BGPV_SF_OUT1, BGPV_SF_OUT2, BGPV_SF_OUT3,
     BGPV_SF_OUT4, BGPV_SF_OUT5, BGPV_SF_OUT6, CLKN_DX, CLKN_SX,
     CLKP_DX, CLKP_SX, 
     /*GNDA_BGPV_MON, GNDA_LBL_MON, GNDA_TO_MON,
     GNDA_WC_BGPV_MON, GNDA_WC_LBL_MON, GNDA_WC_TO_MON, GNDD_BGPV_MON,
     GNDD_LBL_MON, GNDD_TO_MON, GNDD_WC_BGPV_MON, GNDD_WC_LBL_MON,
     GNDD_WC_TO_MON, */
     GND_TOP, LBNL_OUT1_1I, LBNL_OUT1_1O, LBNL_OUT1_2I,
     LBNL_OUT1_2O, LBNL_OUT1_3I, LBNL_OUT1_3O, LBNL_OUT2B_1I,
     LBNL_OUT2B_1O, LBNL_OUT2B_2I, LBNL_OUT2B_2O, LBNL_OUT2B_3I,
     LBNL_OUT2B_3O, LBNL_OUT2_1I, LBNL_OUT2_1O, LBNL_OUT2_2I,
     LBNL_OUT2_2O, LBNL_OUT2_3I, LBNL_OUT2_3O, TO_OE12, TO_OE34,
     TO_OE56, TO_PA1, TO_PA2, TO_PA3, TO_PA4, TO_PA5, TO_PA6, TO_SF_IN,
     TO_SF_OUT, TO_SF_OUT1, TO_SF_OUT2, TO_SF_OUT3, TO_SF_OUT4,
     TO_SF_OUT5, TO_SF_OUT6, 
     /*VDDA_BGPV_MON, VDDA_LBL_MON,
     VDDA_TOP_LBNL, VDDA_TO_MON, VDDA_WC_BGPV_MON, VDDA_WC_LBL_MON,
     VDDA_WC_TO_MON, VDDD_BGPV_MON, VDDD_LBL_MON, VDDD_TO_MON,
     VDDD_WC_BGPV_MON, VDDD_WC_LBL_MON, VDDD_WC_TO_MON,*/
     VDD_CAP_DX, VDD_CAP_SX, VDD_PCAP_DX, VDD_PCAP_SX, VDD_TOP
     /*, VSUB */
     );

inout  BGPV_OE12, BGPV_OE34, BGPV_OE56, BGPV_PA1, BGPV_PA2, BGPV_PA3,
     BGPV_PA4, BGPV_PA5, BGPV_PA6, BGPV_SF_IN, BGPV_SF_OUT,
     BGPV_SF_OUT1, BGPV_SF_OUT2, BGPV_SF_OUT3, BGPV_SF_OUT4,
     BGPV_SF_OUT5, BGPV_SF_OUT6, CLKN_DX, CLKN_SX, CLKP_DX, CLKP_SX,
     
     /*GNDA_BGPV_MON, GNDA_LBL_MON, GNDA_TO_MON, GNDA_WC_BGPV_MON,
     GNDA_WC_LBL_MON, GNDA_WC_TO_MON, GNDD_BGPV_MON, GNDD_LBL_MON,
     GNDD_TO_MON, GNDD_WC_BGPV_MON, GNDD_WC_LBL_MON, GNDD_WC_TO_MON,*/
     
     GND_TOP, LBNL_OUT1_1I, LBNL_OUT1_1O, LBNL_OUT1_2I, LBNL_OUT1_2O,
     LBNL_OUT1_3I, LBNL_OUT1_3O, LBNL_OUT2B_1I, LBNL_OUT2B_1O,
     LBNL_OUT2B_2I, LBNL_OUT2B_2O, LBNL_OUT2B_3I, LBNL_OUT2B_3O,
     LBNL_OUT2_1I, LBNL_OUT2_1O, LBNL_OUT2_2I, LBNL_OUT2_2O,
     LBNL_OUT2_3I, LBNL_OUT2_3O, TO_OE12, TO_OE34, TO_OE56, TO_PA1,
     TO_PA2, TO_PA3, TO_PA4, TO_PA5, TO_PA6, TO_SF_IN, TO_SF_OUT,
     TO_SF_OUT1, TO_SF_OUT2, TO_SF_OUT3, TO_SF_OUT4, TO_SF_OUT5,
     TO_SF_OUT6, 
     
     /*VDDA_BGPV_MON, VDDA_LBL_MON, VDDA_TOP_LBNL,
     VDDA_TO_MON, VDDA_WC_BGPV_MON, VDDA_WC_LBL_MON, VDDA_WC_TO_MON,
     VDDD_BGPV_MON, VDDD_LBL_MON, VDDD_TO_MON, VDDD_WC_BGPV_MON,
     VDDD_WC_LBL_MON, VDDD_WC_TO_MON, */
     
     VDD_CAP_DX, VDD_CAP_SX,
     VDD_PCAP_DX, VDD_PCAP_SX, VDD_TOP; //, VSUB;



endmodule


//-----------------------------------------------------------------------------------------------------
//                                        VLSI Design Laboratory
//                               Istituto Nazionale di Fisica Nucleare (INFN)
//                                   via Giuria 1 10125, Torino, Italy
//-----------------------------------------------------------------------------------------------------
// [Filename]       JTAG_TAP_FSM.sv [RTL]
// [Project]        RD53A pixel ASIC demonstrator
// [Author]         Luca Pacher - pacher@to.infn.it
// [Language]       SystemVerilog 2012 [IEEE Std. 1800-2012]
// [Created]        Jul  4, 2016
// [Modified]       Apr 13, 2017
// [Description]    Fully IEEE Std. 1149.1-2001 compliant JTAG Test Access Port (TAP) FSM controller
//
// [Notes]          Mealy FSM coding style. Hamming protection no more supported/required.
//
// [Status]         devel
//-----------------------------------------------------------------------------------------------------


// Dependencies:
//
// $RTL_DIR/eoc/jtag/TAP_FSM_codes_pkg.sv   **NOTE: package source file included at top-level


`ifndef JTAG_TAP_FSM__SV
`define JTAG_TAP_FSM__SV


`timescale 1ns / 1ps
//`include "timescale.v"


module JTAG_TAP_FSM (

   input  wire TRST,                     // Test Reset (asynchronous, active-low) 
   input  wire TCK,                      // Test Clock
   input  wire TMS,                      // Test Mode Select

   output  logic   SELECT_DR,
   output  logic    SHIFT_DR,            // shift-enable for selected data-register        (right-shift TDI into selected DR shift register)
   output  logic   UPDATE_DR,            // latch-enable for selected data-register        (transfer selected DR shift register data into DR output shadow register)
   output  logic  CAPTURE_DR,            // load-enable  for selected data-register        (load an optional parallel-load into selected DR shift register)
   output  logic    CLOCK_DR,            // shift-enable for boundary-scan registers

   output  logic   SELECT_IR,
   output  logic    SHIFT_IR,            // shift-enable for JTAG instruction-register     (right-shift TDI into IR shift register)
   output  logic   UPDATE_IR,            // latch-enable for JTAG instruction-register     (transfer IR shift register data into IR output shadow register)
   output  logic  CAPTURE_IR,            // load-enable  for JTAG instruction-register     (load an optional parallel-load into IR shift register)

   output  logic  RESET,                 // TAP reset (synchronous with TCK, active-low)
   output  logic  SELECT,                // control signal for TDO_DR/TDO_IR multiplexer
   output  logic  ENABLE                 // control signal for TDO tri-state output buffer

   //output  CLOCK_DR,                   // **NOTE: gated-clocks CLOCK_DR/CLOCK_IR and UPDATE_DR/UPDATE_IR generated from TAP controller not adopted (IEEE Std. 1149.1-2001 broken), they
   //output  CLOCK_IR                    //         are mentioned in RTL just for reference. TCK is propagated to all JTAG clock pins instead

   ) ;


   `ifndef ABSTRACT


   // 4-bit binary-encoded or 15-bit one-hot encoded current/next state types
   import JTAG_TAP_FSM_codes_pkg::* ;

   JTAG_TAP_state STATE ;
   JTAG_TAP_state NEXT_STATE ;


   // internal signals generated by TAP controller (pure combinational outputs)
   logic  SELECT_DR_STATE ;
   logic   SHIFT_DR_STATE ;
   logic  UPDATE_DR_STATE ;
   logic CAPTURE_DR_STATE ;

   logic  SELECT_IR_STATE ;
   logic   SHIFT_IR_STATE ;
   logic  UPDATE_IR_STATE ;
   logic CAPTURE_IR_STATE ;

   logic      RESET_STATE ;
   logic     SELECT_STATE ;

   logic   CLOCK_DR_STATE ;
   logic   CLOCK_IR_STATE ;


   // next_state logic (pure sequential block)
   always_ff @(negedge TRST or posedge TCK) begin

      if( TRST == 1'b0 )
         STATE <= Test_Logic_Reset ;      // active-low asynchronous reset (according to IEEE Std. 1149.1-2001)
      else
         STATE <= NEXT_STATE ;
   end


   // state-transitions and state-outputs table
   // **NOTE: ENABLE = SHIFT_DR | SHIFT_IR

   //-------------------------------------------------------------------------------------------------------------------------------------------
   //                    |                                                  State output ( * = TBC )
   //      TAP state     |----------------------------------------------------------------------------------------------------------------------
   //                    |  CLOCK_DR  CAPTURE_DR  SHIFT_DR  UPDATE_DR  |  CLOCK_IR  CAPTURE_IR  SHIFT_IR  UPDATE_IR   |  RESET  SELECT  ENABLE
   //--------------------|----------------------------------------------------------------------------------------------------------------------
   //  Test Logic Reset  |     0          0           0         0      |      0          0          0          0      |    0      1*      0
   //  Run Test/Idle     |     0          0           0         0      |      0          0          0          0      |    1      1*      0
   //-------------------------------------------------------------------------------------------------------------------------------------------
   //  Select  DR Scan   |     0          0           0         0      |      0          0          0          0      |    1      0       0
   //  Capture DR        |     1          1           0         0      |      0          0          0          0      |    1      0       0
   //  Shift   DR        |     1          0           1         0      |      0          0          0          0      |    1      0       1
   //  Exit1   DR        |     0          0           0         0      |      0          0          0          0      |    1      0       0
   //  Pause   DR        |     0          0           0         0      |      0          0          0          0      |    1      0       0
   //  Exit2   DR        |     0          0           0         0      |      0          0          0          0      |    1      0       0
   //  Update  DR        |     0          0           0         1      |      0          0          0          0      |    1      0       0
   //-------------------------------------------------------------------------------------------------------------------------------------------
   //  Select  IR Scan   |     0          0           0         0      |      0          0          0          0      |    1      1       0
   //  Capture IR        |     0          0           0         0      |      1          1          0          0      |    1      1       0
   //  Shift   IR        |     0          0           0         0      |      1          0          1          0      |    1      1       1
   //  Exit1   IR        |     0          0           0         0      |      0          0          0          0      |    1      1       0
   //  Pause   IR        |     0          0           0         0      |      0          0          0          0      |    1      1       0
   //  Exit2   IR        |     0          0           0         0      |      0          0          0          0      |    1      1       0
   //  Update  IR        |     0          0           0         0      |      0          0          0          1      |    1      1       0
   //-------------------------------------------------------------------------------------------------------------------------------------------

   always_comb begin

       SELECT_DR_STATE = 1'b0 ;
        CLOCK_DR_STATE = 1'b0 ;
      CAPTURE_DR_STATE = 1'b0 ;
        SHIFT_DR_STATE = 1'b0 ;
       UPDATE_DR_STATE = 1'b0 ;

       SELECT_IR_STATE = 1'b0 ;
        CLOCK_IR_STATE = 1'b0 ;
      CAPTURE_IR_STATE = 1'b0 ;
        SHIFT_IR_STATE = 1'b0 ;
       UPDATE_IR_STATE = 1'b0 ;

           RESET_STATE = 1'b0 ;
          SELECT_STATE = 1'b0 ;

      unique case ( STATE )

         //default : NEXT_STATE <= Test_Logic_Reset ;   // catch-all, not required (unique case)


         // Test Logic Reset
         Test_Logic_Reset : begin

             SELECT_DR_STATE = 1'b0 ;
              CLOCK_DR_STATE = 1'b0 ;
            CAPTURE_DR_STATE = 1'b0 ;
              SHIFT_DR_STATE = 1'b0 ;
             UPDATE_DR_STATE = 1'b0 ;

             SELECT_IR_STATE = 1'b0 ;
              CLOCK_IR_STATE = 1'b0 ;
            CAPTURE_IR_STATE = 1'b0 ;
              SHIFT_IR_STATE = 1'b0 ;
             UPDATE_IR_STATE = 1'b0 ;

                 RESET_STATE = 1'b0 ;     // **NOTE: the internal RESET_STATE is active-high, but the re-synched RESET output is inverted, hence active-low    
                SELECT_STATE = 1'b1 ;     // (TBC)


            if( TMS == 1'b1 )
               NEXT_STATE = Test_Logic_Reset ;
            else
               NEXT_STATE = Run_Test_Idle ;
         end

         //______________________________________________________________________
         //


         // Run Test/Idle
         Run_Test_Idle : begin

             SELECT_DR_STATE = 1'b0 ;
              CLOCK_DR_STATE = 1'b0 ;
            CAPTURE_DR_STATE = 1'b0 ;
              SHIFT_DR_STATE = 1'b0 ;
             UPDATE_DR_STATE = 1'b0 ;

             SELECT_IR_STATE = 1'b0 ;
              CLOCK_IR_STATE = 1'b0 ;
            CAPTURE_IR_STATE = 1'b0 ;
              SHIFT_IR_STATE = 1'b0 ;
             UPDATE_IR_STATE = 1'b0 ;

                 RESET_STATE = 1'b1 ;
                SELECT_STATE = 1'b1 ;     // (TBC)


            if( TMS == 1'b1 )
               NEXT_STATE = Select_DR_Scan ;
            else
               NEXT_STATE = Run_Test_Idle ;
         end

         //______________________________________________________________________
         //


         // Select Data Register
         Select_DR_Scan : begin

             SELECT_DR_STATE = 1'b1 ;
              CLOCK_DR_STATE = 1'b0 ;
            CAPTURE_DR_STATE = 1'b0 ;
              SHIFT_DR_STATE = 1'b0 ;
             UPDATE_DR_STATE = 1'b0 ;

             SELECT_IR_STATE = 1'b0 ;
              CLOCK_IR_STATE = 1'b0 ;
            CAPTURE_IR_STATE = 1'b0 ;
              SHIFT_IR_STATE = 1'b0 ;
             UPDATE_IR_STATE = 1'b0 ;

                 RESET_STATE = 1'b1 ;
                SELECT_STATE = 1'b0 ;


            if( TMS == 1'b1 )
               NEXT_STATE = Select_IR_Scan ;
            else
               NEXT_STATE = Capture_DR ;
          end

         //______________________________________________________________________
         //


         // Capture Data Register
         Capture_DR : begin

             SELECT_DR_STATE = 1'b0 ;
              CLOCK_DR_STATE = 1'b1 ;
            CAPTURE_DR_STATE = 1'b1 ;
              SHIFT_DR_STATE = 1'b0 ;
             UPDATE_DR_STATE = 1'b0 ;

             SELECT_IR_STATE = 1'b0 ;
              CLOCK_IR_STATE = 1'b0 ;
            CAPTURE_IR_STATE = 1'b0 ;
              SHIFT_IR_STATE = 1'b0 ;
             UPDATE_IR_STATE = 1'b0 ;

                 RESET_STATE = 1'b1 ;
                SELECT_STATE = 1'b0 ;


            if( TMS == 1'b1 )
               NEXT_STATE = Exit1_DR ;
            else
               NEXT_STATE = Shift_DR ;
         end

         //______________________________________________________________________
         //


         // Shift Data Register
         Shift_DR : begin

             SELECT_DR_STATE = 1'b0 ;
              CLOCK_DR_STATE = 1'b1 ;
            CAPTURE_DR_STATE = 1'b0 ;
              SHIFT_DR_STATE = 1'b1 ;
             UPDATE_DR_STATE = 1'b0 ;

             SELECT_IR_STATE = 1'b0 ;
              CLOCK_IR_STATE = 1'b0 ;
            CAPTURE_IR_STATE = 1'b0 ;
              SHIFT_IR_STATE = 1'b0 ;
             UPDATE_IR_STATE = 1'b0 ;

                 RESET_STATE = 1'b1 ;
                SELECT_STATE = 1'b0 ;


            if( TMS == 1'b1 )
               NEXT_STATE = Exit1_DR ;
            else
               NEXT_STATE = Shift_DR ;
         end

         //______________________________________________________________________
         //


         // Exit1 Data Register (nothing to do)
         Exit1_DR : begin

             SELECT_DR_STATE = 1'b0 ;
              CLOCK_DR_STATE = 1'b0 ;
            CAPTURE_DR_STATE = 1'b0 ;
              SHIFT_DR_STATE = 1'b0 ;
             UPDATE_DR_STATE = 1'b0 ;

             SELECT_IR_STATE = 1'b0 ;
              CLOCK_IR_STATE = 1'b0 ;
            CAPTURE_IR_STATE = 1'b0 ;
              SHIFT_IR_STATE = 1'b0 ;
             UPDATE_IR_STATE = 1'b0 ;

                 RESET_STATE = 1'b1 ;
                SELECT_STATE = 1'b0 ;


            if( TMS == 1'b1 )
               NEXT_STATE = Update_DR ;
            else
               NEXT_STATE = Pause_DR ;
         end

         //______________________________________________________________________
         //


         // Pause Data Register (nothing to do)
         Pause_DR : begin

             SELECT_DR_STATE = 1'b0 ;
              CLOCK_DR_STATE = 1'b0 ;
            CAPTURE_DR_STATE = 1'b0 ;
              SHIFT_DR_STATE = 1'b0 ;
             UPDATE_DR_STATE = 1'b0 ;

             SELECT_IR_STATE = 1'b0 ;
              CLOCK_IR_STATE = 1'b0 ;
            CAPTURE_IR_STATE = 1'b0 ;
              SHIFT_IR_STATE = 1'b0 ;
             UPDATE_IR_STATE = 1'b0 ;

                 RESET_STATE = 1'b1 ;
                SELECT_STATE = 1'b0 ;


            if( TMS == 1'b1 )
               NEXT_STATE = Exit2_DR ;
            else
               NEXT_STATE = Pause_DR ;
         end

         //______________________________________________________________________
         //


         // Exit2 Data Register (nothing to do)
         Exit2_DR : begin

             SELECT_DR_STATE = 1'b0 ;
              CLOCK_DR_STATE = 1'b0 ;
            CAPTURE_DR_STATE = 1'b0 ;
              SHIFT_DR_STATE = 1'b0 ;
             UPDATE_DR_STATE = 1'b0 ;

             SELECT_IR_STATE = 1'b0 ;
              CLOCK_IR_STATE = 1'b0 ;
            CAPTURE_IR_STATE = 1'b0 ;
              SHIFT_IR_STATE = 1'b0 ;
             UPDATE_IR_STATE = 1'b0 ;

                 RESET_STATE = 1'b1 ;
                SELECT_STATE = 1'b0 ;


            if( TMS == 1'b1 )
               NEXT_STATE = Update_DR ;
            else
               NEXT_STATE = Shift_DR ;
         end

         //______________________________________________________________________
         //


         // Update Data Register
         Update_DR : begin

             SELECT_DR_STATE = 1'b0 ;
              CLOCK_DR_STATE = 1'b0 ;
            CAPTURE_DR_STATE = 1'b0 ;
              SHIFT_DR_STATE = 1'b0 ;
             UPDATE_DR_STATE = 1'b1 ;

             SELECT_IR_STATE = 1'b0 ;
              CLOCK_IR_STATE = 1'b0 ;
            CAPTURE_IR_STATE = 1'b0 ;
              SHIFT_IR_STATE = 1'b0 ;
             UPDATE_IR_STATE = 1'b0 ;

                 RESET_STATE = 1'b1 ;
                SELECT_STATE = 1'b0 ;


            if( TMS == 1'b1 )
               NEXT_STATE = Select_DR_Scan ;
            else
               NEXT_STATE = Run_Test_Idle ;
         end

         //______________________________________________________________________
         //


         // Select Instruction Register
         Select_IR_Scan : begin

             SELECT_DR_STATE = 1'b0 ;
              CLOCK_DR_STATE = 1'b0 ;
            CAPTURE_DR_STATE = 1'b0 ;
              SHIFT_DR_STATE = 1'b0 ;
             UPDATE_DR_STATE = 1'b0 ;

             SELECT_IR_STATE = 1'b1 ;
              CLOCK_IR_STATE = 1'b0 ;
            CAPTURE_IR_STATE = 1'b0 ;
              SHIFT_IR_STATE = 1'b0 ;
             UPDATE_IR_STATE = 1'b0 ;

                 RESET_STATE = 1'b1 ;
                SELECT_STATE = 1'b1 ;


            if( TMS == 1'b1 )
               NEXT_STATE = Test_Logic_Reset ;
            else
               NEXT_STATE = Capture_IR ;
         end

         //______________________________________________________________________
         //


         // Capture Instruction Register
         Capture_IR : begin

              CLOCK_DR_STATE = 1'b0 ;
            CAPTURE_DR_STATE = 1'b0 ;
              SHIFT_DR_STATE = 1'b0 ;
             UPDATE_DR_STATE = 1'b0 ;

             SELECT_IR_STATE = 1'b0 ;
              CLOCK_IR_STATE = 1'b1 ;
            CAPTURE_IR_STATE = 1'b1 ;
              SHIFT_IR_STATE = 1'b0 ;
             UPDATE_IR_STATE = 1'b0 ;

                 RESET_STATE = 1'b1 ;
                SELECT_STATE = 1'b1 ;


            if( TMS == 1'b1 )
               NEXT_STATE = Exit1_IR ;
            else
               NEXT_STATE = Shift_IR ;
         end

         //______________________________________________________________________
         //


         // Shift Instruction Register
         Shift_IR : begin

             SELECT_DR_STATE = 1'b0 ;
              CLOCK_DR_STATE = 1'b0 ;
            CAPTURE_DR_STATE = 1'b0 ;
              SHIFT_DR_STATE = 1'b0 ;
             UPDATE_DR_STATE = 1'b0 ;

             SELECT_IR_STATE = 1'b0 ;
              CLOCK_IR_STATE = 1'b1 ;
            CAPTURE_IR_STATE = 1'b0 ;
              SHIFT_IR_STATE = 1'b1 ;
             UPDATE_IR_STATE = 1'b0 ;

                 RESET_STATE = 1'b1 ;
                SELECT_STATE = 1'b1 ;


            if( TMS == 1'b1 )
               NEXT_STATE = Exit1_IR ;
            else
               NEXT_STATE = Shift_IR ;
         end

         //______________________________________________________________________
         //


         // Exit1 Instruction Register (nothing to do, just select IR path)
         Exit1_IR : begin

             SELECT_DR_STATE = 1'b0 ;
              CLOCK_DR_STATE = 1'b0 ;
            CAPTURE_DR_STATE = 1'b0 ;
              SHIFT_DR_STATE = 1'b0 ;
             UPDATE_DR_STATE = 1'b0 ;

             SELECT_IR_STATE = 1'b0 ;
              CLOCK_IR_STATE = 1'b0 ;
            CAPTURE_IR_STATE = 1'b0 ;
              SHIFT_IR_STATE = 1'b0 ;
             UPDATE_IR_STATE = 1'b0 ;

                 RESET_STATE = 1'b1 ;
                SELECT_STATE = 1'b1 ;


            if( TMS == 1'b1 )
               NEXT_STATE = Update_IR ;
            else
               NEXT_STATE = Pause_IR ;
         end

         //______________________________________________________________________
         //


         // Pause Instruction Register (nothing to do, just select IR path)
         Pause_IR : begin

             SELECT_DR_STATE = 1'b0 ;
              CLOCK_DR_STATE = 1'b0 ;
            CAPTURE_DR_STATE = 1'b0 ;
              SHIFT_DR_STATE = 1'b0 ;
             UPDATE_DR_STATE = 1'b0 ;

             SELECT_IR_STATE = 1'b0 ;
              CLOCK_IR_STATE = 1'b0 ;
            CAPTURE_IR_STATE = 1'b0 ;
              SHIFT_IR_STATE = 1'b0 ;
             UPDATE_IR_STATE = 1'b0 ;

                 RESET_STATE = 1'b1 ;
                SELECT_STATE = 1'b1 ;


            if( TMS == 1'b1 )
               NEXT_STATE = Exit2_IR ;
            else
               NEXT_STATE = Pause_IR ;
         end

         //______________________________________________________________________
         //


         // Exit2 Instruction Register (nothing to do, just select IR path)
         Exit2_IR : begin

             SELECT_DR_STATE = 1'b0 ;
              CLOCK_DR_STATE = 1'b0 ;
            CAPTURE_DR_STATE = 1'b0 ;
              SHIFT_DR_STATE = 1'b0 ;
             UPDATE_DR_STATE = 1'b0 ;

             SELECT_IR_STATE = 1'b0 ;
              CLOCK_IR_STATE = 1'b0 ;
            CAPTURE_IR_STATE = 1'b0 ;
              SHIFT_IR_STATE = 1'b0 ;
             UPDATE_IR_STATE = 1'b0 ;

                 RESET_STATE = 1'b1 ;
                SELECT_STATE = 1'b1 ;


            if( TMS == 1'b1 )
               NEXT_STATE = Update_IR ;
            else
               NEXT_STATE = Shift_IR ;
         end

         //______________________________________________________________________
         //


         // Update Instruction Register
         Update_IR : begin

             SELECT_DR_STATE = 1'b0 ;
              CLOCK_DR_STATE = 1'b0 ;
            CAPTURE_DR_STATE = 1'b0 ;
              SHIFT_DR_STATE = 1'b0 ;
             UPDATE_DR_STATE = 1'b0 ;

             SELECT_IR_STATE = 1'b0 ;
              CLOCK_IR_STATE = 1'b0 ;
            CAPTURE_IR_STATE = 1'b0 ;
              SHIFT_IR_STATE = 1'b0 ;
             UPDATE_IR_STATE = 1'b1 ;

                 RESET_STATE = 1'b1 ;
                SELECT_STATE = 1'b1 ;


            if( TMS == 1'b1 )
               NEXT_STATE = Select_DR_Scan ;
            else
               NEXT_STATE = Run_Test_Idle ;
         end

      endcase
   end   // always_comb



   // control signal for TDO tri-state output buffer
   wire   ENABLE_STATE ;
   assign ENABLE_STATE = SHIFT_DR_STATE | SHIFT_IR_STATE ;



   // re-synch all FSM outputs @(negedge TCK) **EXCEPT** UPDATE_DR/UPDATE_IR

   always_ff @(negedge TRST or negedge TCK) begin

      if( TRST == 1'b0 ) begin

          SELECT_DR <= 1'b0 ;
           SHIFT_DR <= 1'b0 ;
         CAPTURE_DR <= 1'b0 ;
           CLOCK_DR <= 1'b0 ;

          SELECT_IR <= 1'b0 ;
           SHIFT_IR <= 1'b0 ;
         CAPTURE_IR <= 1'b0 ;

              RESET <= 1'b0 ;    // **NOTE: TAP reset is also asserted when in Test-Reset-Logic state
             SELECT <= 1'b0 ;
             ENABLE <= 1'b0 ;

      end
      else begin

          SELECT_DR <=   SELECT_DR_STATE ;
           SHIFT_DR <=    SHIFT_DR_STATE ;
         CAPTURE_DR <=  CAPTURE_DR_STATE ;
           CLOCK_DR <=    CLOCK_DR_STATE ;

          SELECT_IR <=   SELECT_IR_STATE ;
           SHIFT_IR <=    SHIFT_IR_STATE ;
         CAPTURE_IR <=  CAPTURE_IR_STATE ;

              RESET <=       RESET_STATE ;
             SELECT <=      SELECT_STATE ;
             ENABLE <=      ENABLE_STATE ;

      end // else
   end  // always_ff



   // re-synch UPDATE_DR/UPDATE_IR FSM outputs @(posedge TCK)

   always_ff @(negedge TRST or posedge TCK) begin

      if( TRST == 1'b0 ) begin

         UPDATE_DR <= 1'b0 ;
         UPDATE_IR <= 1'b0 ;

      end
      else begin

         UPDATE_DR <= UPDATE_DR_STATE ;
         UPDATE_IR <= UPDATE_IR_STATE ;

      end // else
   end   // always_ff

   `endif // ABSTRACT


endmodule : JTAG_TAP_FSM

`endif

